module kyber;
  // this thing should be the top level sytem design but I suck at Verilog programming
  
endmodule