module invntt(
  input clk,
  input set,
  input reset,
  output reg done
); 

endmodule