module cbd2_cal(
  input clk,
  input set,
  input wire [31:0] din,
  output reg [31:0] dout
);

reg [31:0] d;
// TODO: should I make it combinational????
always @(posedge clk) begin
  if(set) begin
    d = (din & 32'h55555555) + ((din >> 1) & 32'h55555555);
    dout =  ((( ((d >> (4*0)) & 'h3) - ((d >> (4*0+2)) & 'h3) ) & 'hf ) << 24 /*0 */ )
          | ((( ((d >> (4*1)) & 'h3) - ((d >> (4*1+2)) & 'h3) ) & 'hf ) << 28 /*4 */ )
          | ((( ((d >> (4*2)) & 'h3) - ((d >> (4*2+2)) & 'h3) ) & 'hf ) << 16 /*8 */ )
          | ((( ((d >> (4*3)) & 'h3) - ((d >> (4*3+2)) & 'h3) ) & 'hf ) << 20 /*12*/ )
          | ((( ((d >> (4*4)) & 'h3) - ((d >> (4*4+2)) & 'h3) ) & 'hf ) <<  8 /*16*/ )
          | ((( ((d >> (4*5)) & 'h3) - ((d >> (4*5+2)) & 'h3) ) & 'hf ) << 12 /*20*/ )
          | ((( ((d >> (4*6)) & 'h3) - ((d >> (4*6+2)) & 'h3) ) & 'hf ) <<  0 /*24*/ )
          | ((( ((d >> (4*7)) & 'h3) - ((d >> (4*7+2)) & 'h3) ) & 'hf ) <<  4 /*28*/ )
          ;
  end
end

endmodule
