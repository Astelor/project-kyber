module cbd(
  input clk,
  
);

endmodule