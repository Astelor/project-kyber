module fifo #(parameter WIDTH = 16)(
  input clk,
  input set,
  input [WIDTH-1:0] wire 
);

endmodule