module invntt(
  input clk,
  input set,
  
); 

endmodule